`timescale 1ns/1ps
`include "KNN_Header.vh"
`include "iob_lib.vh"
 module knn_core
(
  `INPUT(KNN_START_CORE,1),
  `INPUT(KNN_DATA_PT_CORE1,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE2,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE3,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE4,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE5,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE6,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE7,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE8,`WDATA_W),
  `INPUT(KNN_TEST_PT_CORE,`WDATA_W),
  `INPUT(KNN_VALID_CORE,1),
  `INPUT(KNN_SAMPLE_CORE,1),
  `OUTPUT(KNN_VALID_OUT_CORE,1),
 
  `OUTPUT(KN1_OUT_CORE,`WDATA_W),
  `OUTPUT(KN2_OUT_CORE,`WDATA_W),
  `OUTPUT(KN3_OUT_CORE,`WDATA_W),
  `OUTPUT(KN4_OUT_CORE,`WDATA_W),
  `OUTPUT(KN5_OUT_CORE,`WDATA_W),
  `OUTPUT(KN6_OUT_CORE,`WDATA_W),

  `OUTPUT(IN1_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN2_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN3_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN4_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN5_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN6_OUT_CORE,`K_NUM_DATA_PTS_BIT),

  `INPUT(CLK_CORE, 1),
  `INPUT(RST_CORE, 1)

);

`SIGNAL_OUT(KNN_TST_CORE,`WDATA_W)
`SIGNAL_OUT(KNN_DAT_CORE,`WDATA_W)
`SIGNAL_OUT(KNN_ST_CORE,1)

knn_fsm  knn_fsm_inst
(
	//to and from datapath
	.KNN_TEST_PT_O    (KNN_TST_CORE),
	.KNN_DATA_PT_O    (KNN_DAT_CORE),
	.KNN_START_O      (KNN_ST_CORE),
	//to and from KNN top level and KNN core 
	.KNN_START_FSM    (KNN_START_CORE),
	.KNN_DATA_PT_FSM1  (KNN_DATA_PT_CORE1),
	.KNN_DATA_PT_FSM2  (KNN_DATA_PT_CORE2),
	.KNN_DATA_PT_FSM3  (KNN_DATA_PT_CORE3),
	.KNN_DATA_PT_FSM4  (KNN_DATA_PT_CORE4),
	.KNN_DATA_PT_FSM5  (KNN_DATA_PT_CORE5),
	.KNN_DATA_PT_FSM6  (KNN_DATA_PT_CORE6),
	.KNN_DATA_PT_FSM7  (KNN_DATA_PT_CORE7),
	.KNN_DATA_PT_FSM8  (KNN_DATA_PT_CORE8),
	.KNN_TEST_PT_FSM  (KNN_TEST_PT_CORE),
	.KNN_VALID_IN_FSM (KNN_VALID_CORE),
	.KNN_VALID_O      (KNN_VALID_OUT_CORE),
	.clk(CLK_CORE),
	.rst(RST_CORE)
);

knn_datapath knn_datapath_inst
(
	//from fsm
	 .KNN_TEST_PT_DP(KNN_TST_CORE),
	 .KNN_DATA_PT_DP(KNN_DAT_CORE),
	 .KNN_START_DP(KNN_ST_CORE),
	
	//from sw reg
	 .KNN_SAMPLE_DP(KNN_SAMPLE_CORE),
	//to sw reg
	.KN1_OUT(KN1_OUT_CORE),
	.KN2_OUT(KN2_OUT_CORE),
	.KN3_OUT(KN3_OUT_CORE),
	.KN4_OUT(KN4_OUT_CORE),
	.KN5_OUT(KN5_OUT_CORE),
	.KN6_OUT(KN6_OUT_CORE),
	
	.IN1_OUT(IN1_OUT_CORE),
	.IN2_OUT(IN2_OUT_CORE),
	.IN3_OUT(IN3_OUT_CORE),
	.IN4_OUT(IN4_OUT_CORE),
	.IN5_OUT(IN5_OUT_CORE),
	.IN6_OUT(IN6_OUT_CORE),
		
	.clk(CLK_CORE),
	.rst(RST_CORE)
);
		
endmodule 
